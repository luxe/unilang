//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "vend.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w19;    //: /sn:0 {0}(73,522)(117,522){1}
supply0 w4;    //: /sn:0 {0}(480,289)(480,277)(463,277){1}
reg [7:0] w;    //: /sn:0 {0}(#:299,61)(299,146)(362,146)(362,161){1}
reg [7:0] w3;    //: /sn:0 {0}(154,512)(154,483)(#:185,483)(#:185,472){1}
reg w0;    //: /sn:0 {0}(342,381)(205,381)(205,308)(105,308){1}
reg w1;    //: /sn:0 {0}(107,352)(155,352){1}
//: {2}(159,352)(163,352)(163,390)(223,390){3}
//: {4}(157,354)(157,411)(315,411)(315,386)(342,386){5}
reg w8;    //: /sn:0 {0}(543,381)(504,381){1}
//: {2}(500,381)(478,381){3}
//: {4}(502,383)(502,451)(272,451)(272,517)(193,517){5}
supply0 w22;    //: /sn:0 {0}(207,533)(207,527)(193,527){1}
supply0 w12;    //: /sn:0 {0}(534,396)(534,391)(478,391){1}
reg [7:0] w11;    //: /sn:0 {0}(386,161)(386,142)(449,142)(#:449,61){1}
reg w2;    //: /sn:0 {0}(342,391)(319,391)(319,417)(149,417)(149,402){1}
//: {2}(151,400)(223,400){3}
//: {4}(147,400)(111,400){5}
reg [7:0] w10;    //: /sn:0 {0}(#:374,61)(374,161){1}
supply0 [7:0] w9;    //: /sn:0 {0}(#:418,180)(418,154)(398,154)(398,161){1}
supply1 w26;    //: /sn:0 {0}(382,514)(439,514){1}
wire w6;    //: /sn:0 {0}(692,634)(666,634)(666,712)(642,712){1}
wire w7;    //: /sn:0 {0}(309,638)(351,638){1}
//: {2}(355,638)(633,638)(633,611)(692,611){3}
//: {4}(353,636)(353,614){5}
wire w14;    //: /sn:0 {0}(363,386)(402,386){1}
wire [7:0] w16;    //: /sn:0 {0}(#:439,292)(439,376){1}
wire [1:0] w15;    //: /sn:0 {0}(357,177)(258,177)(258,395)(#:229,395){1}
wire w21;    //: /sn:0 {0}(415,277)(400,277){1}
wire [7:0] w20;    //: /sn:0 {0}(#:154,533)(154,558)(287,558)(287,483)(342,483)(342,500){1}
wire [7:0] w23;    //: /sn:0 {0}(#:358,608)(#:358,529){1}
wire w24;    //: /sn:0 {0}(514,686)(606,686)(606,709)(621,709){1}
wire w25;    //: /sn:0 {0}(334,514)(319,514){1}
wire [7:0] w18;    //: /sn:0 {0}(#:439,397)(439,425){1}
//: {2}(#:437,427)(383,427)(383,251)(423,251)(423,263){3}
//: {4}(439,429)(439,487)(374,487)(374,500){5}
wire [7:0] w17;    //: /sn:0 {0}(455,263)(455,237)(380,237)(#:380,190){1}
wire [6:0] w13;    //: /sn:0 {0}(#:493,686)(363,686)(363,614){1}
wire w5;    //: /sn:0 {0}(293,638)(278,638)(278,638)(248,638){1}
//: {2}(244,638)(230,638){3}
//: {4}(246,640)(246,714)(621,714){5}
//: enddecls

  _GGREG8 #(10, 10, 20) g8 (.Q(w18), .D(w16), .EN(w12), .CLR(w8), .CK(w14));   //: @(439,386) /sn:0 /w:[ 0 1 1 3 1 ]
  //: GROUND g4 (w9) @(418,186) /sn:0 /w:[ 0 ]
  //: SWITCH Dime (w1) @(90,352) /w:[ 0 ] /st:0 /dn:0
  //: VDD g13 (w26) @(439,525) /sn:0 /R:3 /w:[ 1 ]
  _GGMUX4x8 #(12, 12) g3 (.I0(w), .I1(w10), .I2(w11), .I3(w9), .S(w15), .Z(w17));   //: @(380,177) /sn:0 /w:[ 1 1 0 1 0 1 ] /ss:0 /do:0
  //: LED Change_Due (w6) @(699,634) /R:3 /w:[ 0 ] /type:0
  //: LED Add_Coin (w7) @(699,611) /R:3 /w:[ 3 ] /type:0
  //: DIP g2 (w11) @(449,51) /sn:0 /w:[ 1 ] /st:25 /dn:0
  //: DIP g1 (w10) @(374,51) /sn:0 /w:[ 0 ] /st:10 /dn:0
  //: LED Vend (w5) @(223,638) /R:1 /w:[ 3 ] /type:0
  _GGNBUF #(2) g16 (.I(w7), .Z(w5));   //: @(303,638) /sn:0 /R:2 /w:[ 0 0 ]
  _GGADD8 #(68, 70, 62, 64) g11 (.A(w18), .B(w17), .S(w16), .CI(w4), .CO(w21));   //: @(439,279) /sn:0 /w:[ 3 0 0 1 0 ]
  //: DIP Price (w3) @(185,462) /w:[ 1 ] /st:100 /dn:0
  //: GROUND g10 (w12) @(534,402) /sn:0 /w:[ 0 ]
  //: joint g19 (w5) @(246, 638) /w:[ 1 -1 2 4 ]
  //: joint g6 (w1) @(157, 352) /w:[ 2 -1 1 4 ]
  //: SWITCH Purchase (w19) @(56,522) /w:[ 0 ] /st:0 /dn:0
  //: joint g9 (w2) @(149, 400) /w:[ 2 -1 4 1 ]
  assign w15 = {w2, w1}; //: CONCAT g7  @(228,395) /sn:0 /w:[ 1 3 3 ] /dr:1 /tp:0 /drp:1
  //: SWITCH Nickel (w0) @(88,308) /w:[ 1 ] /st:0 /dn:0
  //: joint g20 (w7) @(353, 638) /w:[ 2 4 1 -1 ]
  //: DIP Nickel_Amount (w) @(299,51) /sn:0 /w:[ 0 ] /st:5 /dn:0
  assign {w7, w13} = w23; //: CONCAT g15  @(358,609) /sn:0 /R:1 /w:[ 5 1 0 ] /dr:0 /tp:0 /drp:0
  //: SWITCH Quarter (w2) @(94,400) /w:[ 5 ] /st:0 /dn:0
  _GGOR1x7 #(1) g17 (.I0(w13), .Z(w24));   //: @(504,686) /sn:0 /w:[ 0 0 ]
  //: joint g14 (w18) @(439, 427) /w:[ -1 1 2 4 ]
  _GGOR3 #(90) g5 (.I0(w0), .I1(w1), .I2(w2), .Z(w14));   //: @(353,386) /sn:0 /delay:" 90" /w:[ 0 5 0 0 ]
  //: GROUND g24 (w22) @(207,539) /sn:0 /w:[ 0 ]
  _GGREG8 #(10, 10, 20) g21 (.Q(w20), .D(w3), .EN(w22), .CLR(w8), .CK(w19));   //: @(154,522) /sn:0 /w:[ 0 0 1 5 1 ]
  //: SWITCH Reset (w8) @(561,381) /R:2 /w:[ 0 ] /st:1 /dn:0
  //: joint g23 (w8) @(502, 381) /w:[ 1 -1 2 4 ]
  //: GROUND g22 (w4) @(480,295) /sn:0 /w:[ 0 ]
  //: comment g0 @(274,9) /sn:0
  //: /line:"Nickels           Dimes         Quarters"
  //: /end
  _GGADD8 #(70, 72, 62, 64) g12 (.A(~w20), .B(w18), .S(w23), .CI(w26), .CO(w25));   //: @(358,516) /sn:0 /w:[ 1 5 1 0 0 ]
  _GGAND2 #(6) g18 (.I0(w24), .I1(w5), .Z(w6));   //: @(632,712) /sn:0 /w:[ 1 5 1 ]

endmodule
//: /netlistEnd

